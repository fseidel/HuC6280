`default_nettype none

module tb;
  reg clk, reset;
  wire [20:0] AB_21;
  wire [7:0]  DI, DO;
  wire        RE, WE, IRQ, NMI, RDY;
  
  cpu_HuC6280 CPU(.*);
  memory mem(.clk, .re(RE), .we(WE), .addr(AB_21), .dIn(DO), .dOut(DI));

  assign IRQ  = 1'b0;
  assign NMI  = 1'b0;
  assign RDY = 1'b1;

  initial begin
    /*$monitor("AB: %x, DI: %x, PC: %x, State: %s, A: %x, X: %x, Y: %x, S: %x",
             CPU.AB, CPU.DI, CPU.PC, CPU.statename, CPU.A, CPU.X, CPU.Y, CPU.S);*/
    $monitor("AB_21: %x, AB: %x, DI %x, PC: %x, State: %s, MMU_out: %x",
             AB_21, CPU.AB, CPU.DI, CPU.PC, CPU.statename, CPU.MMU_out);
    clk        = 0;
    reset      = 1'b1;
    #10 reset <= 1'b0;
    //#10000 $finish;
    while(CPU.AB != 16'hbeef || ~RE) #10 continue;
    $display("A: %x, X: %x, Y: %x, S: %x",
             CPU.A, CPU.X, CPU.Y, CPU.S);
    #10 $finish;
    //#50000 $finish;
  end

  initial begin
    forever #10 clk = ~clk;
  end

endmodule
